// dummy verilog module for the adjustable oscillator
// TODO How should power and ground be declared?

module osc_adj (
    input vdd,
    input vss,
    input ctrl0,
    input ctrl1,
    output out
);
endmodule
