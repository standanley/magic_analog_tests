magic
tech sky130A
timestamp 1618429821
use test_inverter_adj  test_inverter_adj_0
timestamp 1618341885
transform 1 0 -269 0 1 143
box 260 -145 535 340
<< end >>
