magic
tech sky130A
magscale 1 2
timestamp 1618429821
<< nwell >>
rect 20 420 3460 980
<< metal1 >>
rect 2100 800 2780 860
rect 2880 800 3380 840
rect 2100 760 2140 800
rect 2680 760 2720 800
rect 1680 750 2040 760
rect 1680 690 2000 750
rect 2060 690 2070 750
rect 2180 690 2190 750
rect 2250 690 2260 750
rect 2370 690 2380 750
rect 2440 690 2450 750
rect 2560 690 2570 750
rect 2630 690 2640 750
rect 2750 690 2760 750
rect 2820 690 2830 750
rect 1680 680 2040 690
rect 2100 630 2140 640
rect 1640 550 1680 580
rect 2080 570 2090 630
rect 2150 570 2160 630
rect 2270 570 2280 630
rect 2340 570 2350 630
rect 2460 570 2470 630
rect 2530 570 2540 630
rect 2660 570 2670 630
rect 2730 570 2740 630
rect 1610 530 1680 550
rect 140 340 660 400
rect 740 340 1260 400
rect -20 -40 20 300
rect 1640 50 1680 530
rect 2100 520 2140 570
rect 2680 520 2720 570
rect 2040 460 2720 520
rect 2880 520 2920 800
rect 3060 690 3070 750
rect 3130 690 3140 750
rect 3250 690 3260 750
rect 3320 690 3330 750
rect 2960 570 2970 630
rect 3030 570 3040 630
rect 3160 570 3170 630
rect 3230 570 3240 630
rect 3350 570 3360 630
rect 3420 570 3430 630
rect 2880 480 3280 520
rect 1860 320 1980 380
rect 2060 320 2300 380
rect 2880 360 2920 480
rect 2880 320 3180 360
rect 2284 280 2360 290
rect 1710 220 1720 280
rect 1780 220 1790 280
rect 1900 220 1910 280
rect 1970 220 1980 280
rect 2090 220 2100 280
rect 2160 220 2170 280
rect 2284 220 2370 280
rect 1800 100 1810 160
rect 1870 100 1880 160
rect 2000 100 2010 160
rect 2070 100 2080 160
rect 2190 100 2200 160
rect 2260 100 2270 160
rect 2380 100 2390 160
rect 2450 100 2460 160
rect 2880 60 2920 320
rect 3070 210 3080 270
rect 3140 210 3150 270
rect 2970 100 2980 160
rect 3040 100 3050 160
rect 3160 100 3170 160
rect 3230 100 3240 160
rect 1280 -40 1360 20
rect 1640 10 2390 50
rect 2880 20 3100 60
rect 2880 -40 2920 20
rect -20 -80 2920 -40
<< via1 >>
rect 2000 690 2060 750
rect 2190 690 2250 750
rect 2380 690 2440 750
rect 2570 690 2630 750
rect 2760 690 2820 750
rect 2090 570 2150 630
rect 2280 570 2340 630
rect 2470 570 2530 630
rect 2670 570 2730 630
rect 3070 690 3130 750
rect 3260 690 3320 750
rect 2970 570 3030 630
rect 3170 570 3230 630
rect 3360 570 3420 630
rect 1720 220 1780 280
rect 1910 220 1970 280
rect 2100 220 2160 280
rect 1810 100 1870 160
rect 2010 100 2070 160
rect 2200 100 2260 160
rect 2390 100 2450 160
rect 3080 210 3140 270
rect 2980 100 3040 160
rect 3170 100 3230 160
<< metal2 >>
rect 320 880 1880 940
rect 320 800 380 880
rect 920 800 980 880
rect 1520 800 1580 880
rect 1820 640 1880 880
rect 2000 750 2820 760
rect 2060 690 2190 750
rect 2250 690 2380 750
rect 2440 690 2570 750
rect 2630 690 2760 750
rect 2000 680 2820 690
rect 3070 750 3500 760
rect 3130 690 3260 750
rect 3320 690 3500 750
rect 3070 680 3500 690
rect 1820 630 2150 640
rect 2280 630 2340 640
rect 2470 630 2530 640
rect 2670 630 3420 640
rect 1820 570 2090 630
rect 2150 570 2280 630
rect 2340 570 2470 630
rect 2530 570 2670 630
rect 2730 570 2970 630
rect 3030 570 3170 630
rect 3230 570 3360 630
rect 1820 560 3420 570
rect 1820 290 1880 560
rect 1720 280 2360 290
rect 3460 280 3500 680
rect 1420 170 1480 230
rect 1780 220 1910 280
rect 1970 220 2100 280
rect 2160 220 2360 280
rect 1720 210 2360 220
rect 3080 270 3500 280
rect 3140 210 3500 270
rect 3080 200 3500 210
rect 1420 160 3230 170
rect 1420 100 1810 160
rect 1870 100 2010 160
rect 2070 100 2200 160
rect 2260 100 2390 160
rect 2450 100 2980 160
rect 3040 100 3170 160
rect 1420 90 3230 100
<< metal3 >>
rect 440 560 1740 680
rect 200 160 1480 240
use test_inverter_adj  test_inverter_adj_0
timestamp 1618341885
transform 1 0 -500 0 1 290
box 520 -290 1070 680
use test_inverter_adj  test_inverter_adj_1
timestamp 1618341885
transform 1 0 100 0 1 290
box 520 -290 1070 680
use test_inverter_adj  test_inverter_adj_2
timestamp 1618341885
transform 1 0 700 0 1 290
box 520 -290 1070 680
use sky130_fd_pr__pfet_01v8_RXQGT8  sky130_fd_pr__pfet_01v8_RXQGT8_0
timestamp 1618048189
transform 1 0 2409 0 1 660
box -449 -200 449 200
use sky130_fd_pr__nfet_01v8_PE32AP  sky130_fd_pr__nfet_01v8_PE32AP_0
timestamp 1618046600
transform 1 0 2085 0 1 188
box -365 -188 365 188
use sky130_fd_pr__nfet_01v8_CG72G3  sky130_fd_pr__nfet_01v8_CG72G3_0
timestamp 1618272070
transform 1 0 3105 0 1 188
box -125 -188 125 188
use sky130_fd_pr__pfet_01v8_RX8GT8  sky130_fd_pr__pfet_01v8_RX8GT8_0
timestamp 1618272070
transform 1 0 3197 0 1 660
box -257 -200 257 200
<< labels >>
rlabel metal3 480 600 520 640 1 vdd
port 2 n power bidirectional
rlabel metal3 220 180 260 220 1 vss
port 3 n ground bidirectional
rlabel metal1 1920 320 1980 380 1 ctrl0
port 4 n
rlabel metal1 2160 320 2220 380 1 ctrl1
port 5 n
rlabel metal2 3460 200 3500 760 1 out
port 6 n
<< end >>
