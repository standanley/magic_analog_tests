MACRO test_inverter_adj
  CLASS BLOCK ;
  FOREIGN test_inverter_adj ;
  ORIGIN -2.600 1.450 ;
  SIZE 2.750 BY 4.850 ;
  OBS
      LAYER nwell ;
        RECT 2.600 0.700 4.800 3.400 ;
      LAYER li1 ;
        RECT 3.800 3.080 4.900 3.100 ;
        RECT 3.500 2.900 4.900 3.080 ;
        RECT 3.500 2.620 3.800 2.900 ;
        RECT 2.980 2.435 3.310 2.605 ;
        RECT 4.080 2.435 4.410 2.605 ;
        RECT 4.700 2.220 4.900 2.900 ;
        RECT 2.840 1.180 3.010 2.220 ;
        RECT 3.280 1.180 3.450 2.220 ;
        RECT 3.940 1.180 4.110 2.220 ;
        RECT 4.380 1.900 4.900 2.220 ;
        RECT 4.380 1.180 4.550 1.900 ;
        RECT 2.980 0.795 3.310 0.965 ;
        RECT 4.080 0.795 4.410 0.965 ;
        RECT 3.000 0.230 3.330 0.400 ;
        RECT 2.860 -0.980 3.030 0.060 ;
        RECT 3.300 -0.200 3.470 0.060 ;
        RECT 3.900 -0.200 4.300 -0.120 ;
        RECT 3.300 -0.700 4.300 -0.200 ;
        RECT 3.300 -0.980 3.470 -0.700 ;
        RECT 3.900 -0.780 4.300 -0.700 ;
        RECT 3.000 -1.320 3.330 -1.150 ;
      LAYER mcon ;
        RECT 3.060 2.435 3.230 2.605 ;
        RECT 4.160 2.435 4.330 2.605 ;
        RECT 2.840 1.260 3.010 2.140 ;
        RECT 3.280 1.260 3.450 2.140 ;
        RECT 3.940 1.260 4.110 2.140 ;
        RECT 4.380 1.260 4.550 2.140 ;
        RECT 3.060 0.795 3.230 0.965 ;
        RECT 4.160 0.795 4.330 0.965 ;
        RECT 3.080 0.230 3.250 0.400 ;
        RECT 2.860 -0.900 3.030 -0.020 ;
        RECT 3.300 -0.900 3.470 -0.020 ;
        RECT 3.080 -1.320 3.250 -1.150 ;
      LAYER met1 ;
        RECT 2.950 2.400 3.350 2.700 ;
        RECT 4.050 2.400 4.450 2.700 ;
        RECT 2.810 1.400 3.040 2.200 ;
        RECT 2.600 1.200 3.040 1.400 ;
        RECT 3.250 1.800 3.480 2.200 ;
        RECT 3.910 1.800 4.140 2.200 ;
        RECT 3.250 1.500 4.140 1.800 ;
        RECT 3.250 1.200 3.480 1.500 ;
        RECT 3.910 1.200 4.140 1.500 ;
        RECT 4.350 2.000 4.580 2.200 ;
        RECT 4.350 1.300 5.350 2.000 ;
        RECT 4.350 1.200 4.580 1.300 ;
        RECT 2.600 0.050 2.800 1.200 ;
        RECT 2.950 0.700 3.350 1.000 ;
        RECT 4.050 0.700 4.450 1.000 ;
        RECT 3.000 0.500 3.300 0.700 ;
        RECT 2.950 0.200 3.350 0.500 ;
        RECT 2.600 0.040 3.000 0.050 ;
        RECT 2.600 -0.200 3.060 0.040 ;
        RECT 2.830 -0.960 3.060 -0.200 ;
        RECT 3.270 -0.200 3.500 0.040 ;
        RECT 3.270 -0.700 3.900 -0.200 ;
        RECT 3.270 -0.960 3.500 -0.700 ;
        RECT 2.950 -1.400 3.350 -1.100 ;
      LAYER via ;
        RECT 3.000 2.400 3.300 2.700 ;
        RECT 4.100 2.400 4.400 2.700 ;
        RECT 4.700 1.300 5.300 2.000 ;
        RECT 3.000 0.700 3.300 1.000 ;
        RECT 4.100 0.700 4.400 1.000 ;
        RECT 3.000 0.200 3.300 0.500 ;
        RECT 3.000 -1.400 3.300 -1.100 ;
      LAYER met2 ;
        RECT 3.000 -1.450 3.300 2.750 ;
        RECT 4.100 0.650 4.400 2.750 ;
        RECT 4.700 1.250 5.300 2.050 ;
        RECT 3.500 -0.750 3.900 -0.150 ;
      LAYER via2 ;
        RECT 4.700 1.300 5.300 2.000 ;
        RECT 3.500 -0.700 3.900 -0.200 ;
      LAYER met3 ;
        RECT 4.650 1.275 5.350 2.025 ;
        RECT 3.400 -0.800 4.000 -0.100 ;
  END
END test_inverter_adj
END LIBRARY

