* SPICE3 file created from test_osc_adj.ext - technology: sky130A

.option scale=5000u

.subckt test_osc_adj vdd vss ctrl0 ctrl1 out
X0 out test_inverter_adj_2/in vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X1 out test_inverter_adj_2/in vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X2 vdd test_inverter_adj_2/in out vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X3 vdd test_inverter_adj_2/in out vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X4 test_inverter_adj_2/ctrl ctrl1 vss vss sky130_fd_pr__nfet_01v8 w=200 l=30
X5 vss vdd test_inverter_adj_2/ctrl vss sky130_fd_pr__nfet_01v8 w=200 l=30
X6 test_inverter_adj_2/ctrl ctrl0 vss vss sky130_fd_pr__nfet_01v8 w=200 l=30
X7 vss vdd test_inverter_adj_2/ctrl vss sky130_fd_pr__nfet_01v8 w=200 l=30
X8 test_inverter_adj_2/ctrl ctrl1 vss vss sky130_fd_pr__nfet_01v8 w=200 l=30
X9 vss vdd test_inverter_adj_2/ctrl vss sky130_fd_pr__nfet_01v8 w=200 l=30
X10 vss vdd test_inverter_adj_2/ctrl vss sky130_fd_pr__nfet_01v8 w=200 l=30
X11 vss test_inverter_adj_2/in out vss sky130_fd_pr__nfet_01v8 w=200 l=30
X12 out test_inverter_adj_2/in vss vss sky130_fd_pr__nfet_01v8 w=200 l=30
X13 vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X14 test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X15 vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X16 vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X17 test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X18 vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X19 test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X20 test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X21 vss test_inverter_adj_0/in test_inverter_adj_2/in vss sky130_fd_pr__nfet_01v8 w=200 l=30
X22 test_inverter_adj_0/m1_680_300# test_inverter_adj_0/in test_inverter_adj_2/in vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X23 vdd test_inverter_adj_2/ctrl test_inverter_adj_0/m1_680_300# vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X24 vss test_inverter_adj_1/in test_inverter_adj_0/in vss sky130_fd_pr__nfet_01v8 w=200 l=30
X25 test_inverter_adj_1/m1_680_300# test_inverter_adj_1/in test_inverter_adj_0/in vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X26 vdd test_inverter_adj_2/ctrl test_inverter_adj_1/m1_680_300# vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X27 vss test_inverter_adj_2/in test_inverter_adj_1/in vss sky130_fd_pr__nfet_01v8 w=200 l=30
X28 test_inverter_adj_2/m1_680_300# test_inverter_adj_2/in test_inverter_adj_1/in vdd sky130_fd_pr__pfet_01v8 w=200 l=30
X29 vdd test_inverter_adj_2/ctrl test_inverter_adj_2/m1_680_300# vdd sky130_fd_pr__pfet_01v8 w=200 l=30
C0 test_inverter_adj_2/ctrl vdd 9.13fF
C1 ctrl0 ctrl1 0.07fF
C2 test_inverter_adj_2/ctrl test_inverter_adj_2/in 0.67fF
C3 test_inverter_adj_2/in vdd 1.78fF
C4 test_inverter_adj_1/in test_inverter_adj_1/m1_680_300# 0.39fF
C5 test_inverter_adj_1/in test_inverter_adj_2/m1_680_300# 0.41fF
C6 out test_inverter_adj_2/ctrl 0.08fF
C7 out vdd 2.62fF
C8 test_inverter_adj_0/m1_680_300# test_inverter_adj_0/in 0.39fF
C9 test_inverter_adj_1/in test_inverter_adj_0/in 0.84fF
C10 ctrl0 test_inverter_adj_2/ctrl 0.23fF
C11 ctrl0 vdd 0.10fF
C12 out test_inverter_adj_2/in 0.92fF
C13 ctrl0 test_inverter_adj_2/in 0.01fF
C14 test_inverter_adj_0/m1_680_300# test_inverter_adj_2/ctrl 0.29fF
C15 test_inverter_adj_0/m1_680_300# vdd 0.43fF
C16 test_inverter_adj_1/in test_inverter_adj_2/ctrl 0.55fF
C17 test_inverter_adj_1/in vdd 0.68fF
C18 test_inverter_adj_0/m1_680_300# test_inverter_adj_2/in 0.41fF
C19 test_inverter_adj_1/in test_inverter_adj_2/in 1.00fF
C20 test_inverter_adj_0/in test_inverter_adj_1/m1_680_300# 0.41fF
C21 test_inverter_adj_2/ctrl ctrl1 0.41fF
C22 ctrl1 vdd 0.16fF
C23 test_inverter_adj_1/m1_680_300# test_inverter_adj_2/ctrl 0.29fF
C24 test_inverter_adj_1/m1_680_300# vdd 0.75fF
C25 test_inverter_adj_2/in ctrl1 0.03fF
C26 test_inverter_adj_2/ctrl test_inverter_adj_2/m1_680_300# 0.29fF
C27 test_inverter_adj_2/m1_680_300# vdd 0.78fF
C28 test_inverter_adj_0/in test_inverter_adj_2/ctrl 0.36fF
C29 test_inverter_adj_0/in vdd 0.42fF
C30 test_inverter_adj_2/m1_680_300# test_inverter_adj_2/in 0.30fF
C31 test_inverter_adj_0/in test_inverter_adj_2/in 1.04fF
C32 test_inverter_adj_2/m1_680_300# vss 0.17fF
C33 test_inverter_adj_1/m1_680_300# vss 0.17fF
C34 test_inverter_adj_1/in vss 2.27fF
C35 vdd vss 11.76fF
C36 test_inverter_adj_0/m1_680_300# vss 0.17fF
C37 test_inverter_adj_2/in vss 4.60fF
C38 test_inverter_adj_0/in vss 2.16fF
C39 test_inverter_adj_2/ctrl vss 6.78fF
C40 out vss 1.72fF
C41 ctrl1 vss 0.52fF
C42 ctrl0 vss 0.24fF
.ends
