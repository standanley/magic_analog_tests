magic
tech sky130A
magscale 1 2
timestamp 1618048189
<< error_p >>
rect -269 181 -211 187
rect -77 181 -19 187
rect 115 181 173 187
rect 307 181 365 187
rect -269 147 -257 181
rect -77 147 -65 181
rect 115 147 127 181
rect 307 147 319 181
rect -269 141 -211 147
rect -77 141 -19 147
rect 115 141 173 147
rect 307 141 365 147
rect -365 -147 -307 -141
rect -173 -147 -115 -141
rect 19 -147 77 -141
rect 211 -147 269 -141
rect -365 -181 -353 -147
rect -173 -181 -161 -147
rect 19 -181 31 -147
rect 211 -181 223 -147
rect -365 -187 -307 -181
rect -173 -187 -115 -181
rect 19 -187 77 -181
rect 211 -187 269 -181
<< nwell >>
rect -353 162 449 200
rect -449 -162 449 162
rect -449 -200 353 -162
<< pmos >>
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
<< pdiff >>
rect -413 88 -351 100
rect -413 -88 -401 88
rect -367 -88 -351 88
rect -413 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 413 100
rect 351 -88 367 88
rect 401 -88 413 88
rect 351 -100 413 -88
<< pdiffc >>
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
<< poly >>
rect -273 181 -207 197
rect -273 147 -257 181
rect -223 147 -207 181
rect -273 131 -207 147
rect -81 181 -15 197
rect -81 147 -65 181
rect -31 147 -15 181
rect -81 131 -15 147
rect 111 181 177 197
rect 111 147 127 181
rect 161 147 177 181
rect 111 131 177 147
rect 303 181 369 197
rect 303 147 319 181
rect 353 147 369 181
rect 303 131 369 147
rect -351 100 -321 126
rect -255 100 -225 131
rect -159 100 -129 126
rect -63 100 -33 131
rect 33 100 63 126
rect 129 100 159 131
rect 225 100 255 126
rect 321 100 351 131
rect -351 -131 -321 -100
rect -255 -126 -225 -100
rect -159 -131 -129 -100
rect -63 -126 -33 -100
rect 33 -131 63 -100
rect 129 -126 159 -100
rect 225 -131 255 -100
rect 321 -126 351 -100
rect -369 -147 -303 -131
rect -369 -181 -353 -147
rect -319 -181 -303 -147
rect -369 -197 -303 -181
rect -177 -147 -111 -131
rect -177 -181 -161 -147
rect -127 -181 -111 -147
rect -177 -197 -111 -181
rect 15 -147 81 -131
rect 15 -181 31 -147
rect 65 -181 81 -147
rect 15 -197 81 -181
rect 207 -147 273 -131
rect 207 -181 223 -147
rect 257 -181 273 -147
rect 207 -197 273 -181
<< polycont >>
rect -257 147 -223 181
rect -65 147 -31 181
rect 127 147 161 181
rect 319 147 353 181
rect -353 -181 -319 -147
rect -161 -181 -127 -147
rect 31 -181 65 -147
rect 223 -181 257 -147
<< locali >>
rect -273 147 -257 181
rect -223 147 -207 181
rect -81 147 -65 181
rect -31 147 -15 181
rect 111 147 127 181
rect 161 147 177 181
rect 303 147 319 181
rect 353 147 369 181
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect -369 -181 -353 -147
rect -319 -181 -303 -147
rect -177 -181 -161 -147
rect -127 -181 -111 -147
rect 15 -181 31 -147
rect 65 -181 81 -147
rect 207 -181 223 -147
rect 257 -181 273 -147
<< viali >>
rect -257 147 -223 181
rect -65 147 -31 181
rect 127 147 161 181
rect 319 147 353 181
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect -353 -181 -319 -147
rect -161 -181 -127 -147
rect 31 -181 65 -147
rect 223 -181 257 -147
<< metal1 >>
rect -269 181 -211 187
rect -269 147 -257 181
rect -223 147 -211 181
rect -269 141 -211 147
rect -77 181 -19 187
rect -77 147 -65 181
rect -31 147 -19 181
rect -77 141 -19 147
rect 115 181 173 187
rect 115 147 127 181
rect 161 147 173 181
rect 115 141 173 147
rect 307 181 365 187
rect 307 147 319 181
rect 353 147 365 181
rect 307 141 365 147
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect -365 -147 -307 -141
rect -365 -181 -353 -147
rect -319 -181 -307 -147
rect -365 -187 -307 -181
rect -173 -147 -115 -141
rect -173 -181 -161 -147
rect -127 -181 -115 -147
rect -173 -187 -115 -181
rect 19 -147 77 -141
rect 19 -181 31 -147
rect 65 -181 77 -147
rect 19 -187 77 -181
rect 211 -147 269 -141
rect 211 -181 223 -147
rect 257 -181 269 -147
rect 211 -187 269 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
