magic
tech sky130A
magscale 1 2
timestamp 1618048189
<< error_p >>
rect -29 1707 29 1713
rect -29 1673 -17 1707
rect -29 1667 29 1673
rect -109 1326 109 1544
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect -29 1231 29 1237
rect -109 890 109 1108
rect -29 835 29 841
rect -29 801 -17 835
rect -29 795 29 801
rect -109 454 109 672
rect -29 399 29 405
rect -29 365 -17 399
rect -29 359 29 365
rect -109 18 109 236
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -109 -418 109 -200
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect -29 -513 29 -507
rect -109 -854 109 -636
rect -29 -909 29 -903
rect -29 -943 -17 -909
rect -29 -949 29 -943
rect -109 -1290 109 -1072
rect -29 -1345 29 -1339
rect -29 -1379 -17 -1345
rect -29 -1385 29 -1379
rect -29 -1673 29 -1667
rect -29 -1707 -17 -1673
rect -29 -1713 29 -1707
<< nwell >>
rect -109 1326 109 1726
rect -109 890 109 1290
rect -109 454 109 854
rect -109 18 109 418
rect -109 -418 109 -18
rect -109 -854 109 -454
rect -109 -1290 109 -890
rect -109 -1726 109 -1326
<< pmos >>
rect -15 1426 15 1626
rect -15 990 15 1190
rect -15 554 15 754
rect -15 118 15 318
rect -15 -318 15 -118
rect -15 -754 15 -554
rect -15 -1190 15 -990
rect -15 -1626 15 -1426
<< pdiff >>
rect -73 1614 -15 1626
rect -73 1438 -61 1614
rect -27 1438 -15 1614
rect -73 1426 -15 1438
rect 15 1614 73 1626
rect 15 1438 27 1614
rect 61 1438 73 1614
rect 15 1426 73 1438
rect -73 1178 -15 1190
rect -73 1002 -61 1178
rect -27 1002 -15 1178
rect -73 990 -15 1002
rect 15 1178 73 1190
rect 15 1002 27 1178
rect 61 1002 73 1178
rect 15 990 73 1002
rect -73 742 -15 754
rect -73 566 -61 742
rect -27 566 -15 742
rect -73 554 -15 566
rect 15 742 73 754
rect 15 566 27 742
rect 61 566 73 742
rect 15 554 73 566
rect -73 306 -15 318
rect -73 130 -61 306
rect -27 130 -15 306
rect -73 118 -15 130
rect 15 306 73 318
rect 15 130 27 306
rect 61 130 73 306
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -306 -61 -130
rect -27 -306 -15 -130
rect -73 -318 -15 -306
rect 15 -130 73 -118
rect 15 -306 27 -130
rect 61 -306 73 -130
rect 15 -318 73 -306
rect -73 -566 -15 -554
rect -73 -742 -61 -566
rect -27 -742 -15 -566
rect -73 -754 -15 -742
rect 15 -566 73 -554
rect 15 -742 27 -566
rect 61 -742 73 -566
rect 15 -754 73 -742
rect -73 -1002 -15 -990
rect -73 -1178 -61 -1002
rect -27 -1178 -15 -1002
rect -73 -1190 -15 -1178
rect 15 -1002 73 -990
rect 15 -1178 27 -1002
rect 61 -1178 73 -1002
rect 15 -1190 73 -1178
rect -73 -1438 -15 -1426
rect -73 -1614 -61 -1438
rect -27 -1614 -15 -1438
rect -73 -1626 -15 -1614
rect 15 -1438 73 -1426
rect 15 -1614 27 -1438
rect 61 -1614 73 -1438
rect 15 -1626 73 -1614
<< pdiffc >>
rect -61 1438 -27 1614
rect 27 1438 61 1614
rect -61 1002 -27 1178
rect 27 1002 61 1178
rect -61 566 -27 742
rect 27 566 61 742
rect -61 130 -27 306
rect 27 130 61 306
rect -61 -306 -27 -130
rect 27 -306 61 -130
rect -61 -742 -27 -566
rect 27 -742 61 -566
rect -61 -1178 -27 -1002
rect 27 -1178 61 -1002
rect -61 -1614 -27 -1438
rect 27 -1614 61 -1438
<< poly >>
rect -33 1707 33 1723
rect -33 1673 -17 1707
rect 17 1673 33 1707
rect -33 1657 33 1673
rect -15 1626 15 1657
rect -15 1395 15 1426
rect -33 1379 33 1395
rect -33 1345 -17 1379
rect 17 1345 33 1379
rect -33 1329 33 1345
rect -33 1271 33 1287
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -33 1221 33 1237
rect -15 1190 15 1221
rect -15 959 15 990
rect -33 943 33 959
rect -33 909 -17 943
rect 17 909 33 943
rect -33 893 33 909
rect -33 835 33 851
rect -33 801 -17 835
rect 17 801 33 835
rect -33 785 33 801
rect -15 754 15 785
rect -15 523 15 554
rect -33 507 33 523
rect -33 473 -17 507
rect 17 473 33 507
rect -33 457 33 473
rect -33 399 33 415
rect -33 365 -17 399
rect 17 365 33 399
rect -33 349 33 365
rect -15 318 15 349
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -349 15 -318
rect -33 -365 33 -349
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -415 33 -399
rect -33 -473 33 -457
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -33 -523 33 -507
rect -15 -554 15 -523
rect -15 -785 15 -754
rect -33 -801 33 -785
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -33 -851 33 -835
rect -33 -909 33 -893
rect -33 -943 -17 -909
rect 17 -943 33 -909
rect -33 -959 33 -943
rect -15 -990 15 -959
rect -15 -1221 15 -1190
rect -33 -1237 33 -1221
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -33 -1287 33 -1271
rect -33 -1345 33 -1329
rect -33 -1379 -17 -1345
rect 17 -1379 33 -1345
rect -33 -1395 33 -1379
rect -15 -1426 15 -1395
rect -15 -1657 15 -1626
rect -33 -1673 33 -1657
rect -33 -1707 -17 -1673
rect 17 -1707 33 -1673
rect -33 -1723 33 -1707
<< polycont >>
rect -17 1673 17 1707
rect -17 1345 17 1379
rect -17 1237 17 1271
rect -17 909 17 943
rect -17 801 17 835
rect -17 473 17 507
rect -17 365 17 399
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -17 -835 17 -801
rect -17 -943 17 -909
rect -17 -1271 17 -1237
rect -17 -1379 17 -1345
rect -17 -1707 17 -1673
<< locali >>
rect -33 1673 -17 1707
rect 17 1673 33 1707
rect -61 1614 -27 1630
rect -61 1422 -27 1438
rect 27 1614 61 1630
rect 27 1422 61 1438
rect -33 1345 -17 1379
rect 17 1345 33 1379
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -61 1178 -27 1194
rect -61 986 -27 1002
rect 27 1178 61 1194
rect 27 986 61 1002
rect -33 909 -17 943
rect 17 909 33 943
rect -33 801 -17 835
rect 17 801 33 835
rect -61 742 -27 758
rect -61 550 -27 566
rect 27 742 61 758
rect 27 550 61 566
rect -33 473 -17 507
rect 17 473 33 507
rect -33 365 -17 399
rect 17 365 33 399
rect -61 306 -27 322
rect -61 114 -27 130
rect 27 306 61 322
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -322 -27 -306
rect 27 -130 61 -114
rect 27 -322 61 -306
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -61 -566 -27 -550
rect -61 -758 -27 -742
rect 27 -566 61 -550
rect 27 -758 61 -742
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -33 -943 -17 -909
rect 17 -943 33 -909
rect -61 -1002 -27 -986
rect -61 -1194 -27 -1178
rect 27 -1002 61 -986
rect 27 -1194 61 -1178
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -33 -1379 -17 -1345
rect 17 -1379 33 -1345
rect -61 -1438 -27 -1422
rect -61 -1630 -27 -1614
rect 27 -1438 61 -1422
rect 27 -1630 61 -1614
rect -33 -1707 -17 -1673
rect 17 -1707 33 -1673
<< viali >>
rect -17 1673 17 1707
rect -61 1438 -27 1614
rect 27 1438 61 1614
rect -17 1345 17 1379
rect -17 1237 17 1271
rect -61 1002 -27 1178
rect 27 1002 61 1178
rect -17 909 17 943
rect -17 801 17 835
rect -61 566 -27 742
rect 27 566 61 742
rect -17 473 17 507
rect -17 365 17 399
rect -61 130 -27 306
rect 27 130 61 306
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -306 -27 -130
rect 27 -306 61 -130
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -61 -742 -27 -566
rect 27 -742 61 -566
rect -17 -835 17 -801
rect -17 -943 17 -909
rect -61 -1178 -27 -1002
rect 27 -1178 61 -1002
rect -17 -1271 17 -1237
rect -17 -1379 17 -1345
rect -61 -1614 -27 -1438
rect 27 -1614 61 -1438
rect -17 -1707 17 -1673
<< metal1 >>
rect -29 1707 29 1713
rect -29 1673 -17 1707
rect 17 1673 29 1707
rect -29 1667 29 1673
rect -67 1614 -21 1626
rect -67 1438 -61 1614
rect -27 1438 -21 1614
rect -67 1426 -21 1438
rect 21 1614 67 1626
rect 21 1438 27 1614
rect 61 1438 67 1614
rect 21 1426 67 1438
rect -29 1379 29 1385
rect -29 1345 -17 1379
rect 17 1345 29 1379
rect -29 1339 29 1345
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect 17 1237 29 1271
rect -29 1231 29 1237
rect -67 1178 -21 1190
rect -67 1002 -61 1178
rect -27 1002 -21 1178
rect -67 990 -21 1002
rect 21 1178 67 1190
rect 21 1002 27 1178
rect 61 1002 67 1178
rect 21 990 67 1002
rect -29 943 29 949
rect -29 909 -17 943
rect 17 909 29 943
rect -29 903 29 909
rect -29 835 29 841
rect -29 801 -17 835
rect 17 801 29 835
rect -29 795 29 801
rect -67 742 -21 754
rect -67 566 -61 742
rect -27 566 -21 742
rect -67 554 -21 566
rect 21 742 67 754
rect 21 566 27 742
rect 61 566 67 742
rect 21 554 67 566
rect -29 507 29 513
rect -29 473 -17 507
rect 17 473 29 507
rect -29 467 29 473
rect -29 399 29 405
rect -29 365 -17 399
rect 17 365 29 399
rect -29 359 29 365
rect -67 306 -21 318
rect -67 130 -61 306
rect -27 130 -21 306
rect -67 118 -21 130
rect 21 306 67 318
rect 21 130 27 306
rect 61 130 67 306
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -306 -61 -130
rect -27 -306 -21 -130
rect -67 -318 -21 -306
rect 21 -130 67 -118
rect 21 -306 27 -130
rect 61 -306 67 -130
rect 21 -318 67 -306
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect 17 -399 29 -365
rect -29 -405 29 -399
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect 17 -507 29 -473
rect -29 -513 29 -507
rect -67 -566 -21 -554
rect -67 -742 -61 -566
rect -27 -742 -21 -566
rect -67 -754 -21 -742
rect 21 -566 67 -554
rect 21 -742 27 -566
rect 61 -742 67 -566
rect 21 -754 67 -742
rect -29 -801 29 -795
rect -29 -835 -17 -801
rect 17 -835 29 -801
rect -29 -841 29 -835
rect -29 -909 29 -903
rect -29 -943 -17 -909
rect 17 -943 29 -909
rect -29 -949 29 -943
rect -67 -1002 -21 -990
rect -67 -1178 -61 -1002
rect -27 -1178 -21 -1002
rect -67 -1190 -21 -1178
rect 21 -1002 67 -990
rect 21 -1178 27 -1002
rect 61 -1178 67 -1002
rect 21 -1190 67 -1178
rect -29 -1237 29 -1231
rect -29 -1271 -17 -1237
rect 17 -1271 29 -1237
rect -29 -1277 29 -1271
rect -29 -1345 29 -1339
rect -29 -1379 -17 -1345
rect 17 -1379 29 -1345
rect -29 -1385 29 -1379
rect -67 -1438 -21 -1426
rect -67 -1614 -61 -1438
rect -27 -1614 -21 -1438
rect -67 -1626 -21 -1614
rect 21 -1438 67 -1426
rect 21 -1614 27 -1438
rect 61 -1614 67 -1438
rect 21 -1626 67 -1614
rect -29 -1673 29 -1667
rect -29 -1707 -17 -1673
rect 17 -1707 29 -1673
rect -29 -1713 29 -1707
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 0.15 m 8 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
