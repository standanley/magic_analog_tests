* NGSPICE file created from test_osc_adj.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_RX8GT8 VSUBS a_n33_n100# w_n257_n200# a_n177_n197#
+ a_n81_131# a_15_n197# a_63_n100# a_n221_n100# a_n129_n100# a_111_131# a_159_n100#
X0 a_159_n100# a_111_131# a_63_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_n33_n100# a_n81_131# a_n129_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_n129_n100# a_n177_n197# a_n221_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 a_63_n100# a_15_n197# a_n33_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
C0 a_111_131# a_63_n100# 0.01fF
C1 a_n81_131# a_n177_n197# 0.02fF
C2 a_159_n100# a_n33_n100# 0.11fF
C3 a_n221_n100# a_n33_n100# 0.11fF
C4 a_15_n197# a_n33_n100# 0.01fF
C5 w_n257_n200# a_n33_n100# 0.00fF
C6 a_159_n100# a_n129_n100# 0.06fF
C7 a_n221_n100# a_n129_n100# 0.29fF
C8 a_63_n100# a_n33_n100# 0.29fF
C9 a_n129_n100# w_n257_n200# 0.00fF
C10 a_n221_n100# a_n177_n197# 0.01fF
C11 a_15_n197# a_n177_n197# 0.04fF
C12 a_15_n197# a_n81_131# 0.02fF
C13 a_n129_n100# a_63_n100# 0.11fF
C14 a_159_n100# a_n221_n100# 0.05fF
C15 a_159_n100# w_n257_n200# 0.00fF
C16 a_n221_n100# w_n257_n200# 0.00fF
C17 a_159_n100# a_63_n100# 0.29fF
C18 a_n221_n100# a_63_n100# 0.06fF
C19 a_15_n197# a_63_n100# 0.01fF
C20 w_n257_n200# a_63_n100# 0.00fF
C21 a_111_131# a_n177_n197# 0.00fF
C22 a_n81_131# a_111_131# 0.04fF
C23 a_n129_n100# a_n33_n100# 0.29fF
C24 a_159_n100# a_111_131# 0.01fF
C25 a_n81_131# a_n33_n100# 0.01fF
C26 a_15_n197# a_111_131# 0.02fF
C27 a_n129_n100# a_n177_n197# 0.01fF
C28 a_n129_n100# a_n81_131# 0.01fF
C29 a_159_n100# VSUBS 0.03fF
C30 a_63_n100# VSUBS 0.03fF
C31 a_n33_n100# VSUBS 0.03fF
C32 a_n129_n100# VSUBS 0.03fF
C33 a_n221_n100# VSUBS 0.03fF
C34 a_15_n197# VSUBS 0.12fF
C35 a_n177_n197# VSUBS 0.12fF
C36 a_111_131# VSUBS 0.12fF
C37 a_n81_131# VSUBS 0.12fF
C38 w_n257_n200# VSUBS 0.59fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PE32AP VSUBS a_63_n188# a_n129_n188# a_n81_n100# a_255_n188#
+ a_n273_n100# a_n225_122# a_111_n100# a_n177_n100# a_n33_122# a_15_n100# a_159_122#
+ a_303_n100# a_n321_n188# a_207_n100# a_n365_n100#
X0 a_15_n100# a_n33_122# a_n81_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X1 a_n273_n100# a_n321_n188# a_n365_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X2 a_n177_n100# a_n225_122# a_n273_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X3 a_303_n100# a_255_n188# a_207_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X4 a_207_n100# a_159_122# a_111_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X5 a_n81_n100# a_n129_n188# a_n177_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X6 a_111_n100# a_63_n188# a_15_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
C0 a_n81_n100# a_n365_n100# 0.06fF
C1 a_n81_n100# a_n33_122# 0.01fF
C2 a_n81_n100# a_303_n100# 0.05fF
C3 a_n81_n100# a_n273_n100# 0.11fF
C4 a_15_n100# a_n177_n100# 0.11fF
C5 a_159_122# a_255_n188# 0.02fF
C6 a_63_n188# a_n225_122# 0.00fF
C7 a_63_n188# a_159_122# 0.02fF
C8 a_207_n100# a_255_n188# 0.01fF
C9 a_n177_n100# a_n81_n100# 0.29fF
C10 a_n33_122# a_n225_122# 0.04fF
C11 a_159_122# a_n33_122# 0.04fF
C12 a_n273_n100# a_n225_122# 0.01fF
C13 a_15_n100# a_n81_n100# 0.29fF
C14 a_303_n100# a_207_n100# 0.29fF
C15 a_63_n188# a_n321_n188# 0.02fF
C16 a_n129_n188# a_255_n188# 0.02fF
C17 a_n129_n188# a_63_n188# 0.04fF
C18 a_n177_n100# a_n225_122# 0.01fF
C19 a_n365_n100# a_n321_n188# 0.01fF
C20 a_n33_122# a_n321_n188# 0.00fF
C21 a_63_n188# a_111_n100# 0.01fF
C22 a_n177_n100# a_207_n100# 0.05fF
C23 a_n273_n100# a_n321_n188# 0.01fF
C24 a_n129_n188# a_n33_122# 0.02fF
C25 a_15_n100# a_207_n100# 0.11fF
C26 a_303_n100# a_111_n100# 0.11fF
C27 a_111_n100# a_n273_n100# 0.05fF
C28 a_n129_n188# a_n177_n100# 0.01fF
C29 a_n81_n100# a_207_n100# 0.06fF
C30 a_n177_n100# a_111_n100# 0.06fF
C31 a_63_n188# a_255_n188# 0.04fF
C32 a_159_122# a_n225_122# 0.02fF
C33 a_15_n100# a_111_n100# 0.29fF
C34 a_159_122# a_207_n100# 0.01fF
C35 a_n33_122# a_255_n188# 0.00fF
C36 a_63_n188# a_n33_122# 0.02fF
C37 a_n129_n188# a_n81_n100# 0.01fF
C38 a_303_n100# a_255_n188# 0.01fF
C39 a_n81_n100# a_111_n100# 0.11fF
C40 a_n365_n100# a_n273_n100# 0.29fF
C41 a_n225_122# a_n321_n188# 0.02fF
C42 a_n129_n188# a_n225_122# 0.02fF
C43 a_n129_n188# a_159_122# 0.00fF
C44 a_159_122# a_111_n100# 0.01fF
C45 a_15_n100# a_63_n188# 0.01fF
C46 a_n177_n100# a_n365_n100# 0.11fF
C47 a_n177_n100# a_n273_n100# 0.29fF
C48 a_111_n100# a_207_n100# 0.29fF
C49 a_15_n100# a_n365_n100# 0.05fF
C50 a_15_n100# a_n33_122# 0.01fF
C51 a_15_n100# a_303_n100# 0.06fF
C52 a_15_n100# a_n273_n100# 0.06fF
C53 a_n129_n188# a_n321_n188# 0.04fF
C54 a_303_n100# VSUBS 0.03fF
C55 a_207_n100# VSUBS 0.03fF
C56 a_111_n100# VSUBS 0.03fF
C57 a_15_n100# VSUBS 0.03fF
C58 a_n81_n100# VSUBS 0.03fF
C59 a_n177_n100# VSUBS 0.03fF
C60 a_n273_n100# VSUBS 0.03fF
C61 a_n365_n100# VSUBS 0.03fF
C62 a_255_n188# VSUBS 0.12fF
C63 a_63_n188# VSUBS 0.12fF
C64 a_159_122# VSUBS 0.12fF
C65 a_n129_n188# VSUBS 0.12fF
C66 a_n33_122# VSUBS 0.12fF
C67 a_n321_n188# VSUBS 0.12fF
C68 a_n225_122# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CG72G3 VSUBS a_n33_n100# a_63_n100# a_n81_n188# a_n125_n100#
+ a_15_122#
X0 a_63_n100# a_15_122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n188# a_n125_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
C0 a_n125_n100# a_n81_n188# 0.01fF
C1 a_n33_n100# a_15_122# 0.01fF
C2 a_n33_n100# a_63_n100# 0.29fF
C3 a_15_122# a_63_n100# 0.01fF
C4 a_n33_n100# a_n81_n188# 0.01fF
C5 a_n81_n188# a_15_122# 0.02fF
C6 a_n33_n100# a_n125_n100# 0.29fF
C7 a_n125_n100# a_63_n100# 0.11fF
C8 a_63_n100# VSUBS 0.03fF
C9 a_n33_n100# VSUBS 0.03fF
C10 a_n125_n100# VSUBS 0.03fF
C11 a_n81_n188# VSUBS 0.12fF
C12 a_15_122# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_RXQGT8 VSUBS a_n33_n100# a_n321_n100# a_n273_131#
+ a_n177_n197# a_n81_131# a_15_n197# a_n225_n100# w_n449_n200# a_63_n100# a_n129_n100#
+ a_303_131# a_n369_n197# a_351_n100# a_207_n197# a_255_n100# a_111_131# a_n413_n100#
+ a_159_n100#
X0 a_351_n100# a_303_131# a_255_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_255_n100# a_207_n197# a_159_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_159_n100# a_111_131# a_63_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 a_n33_n100# a_n81_131# a_n129_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 a_n321_n100# a_n369_n197# a_n413_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_n225_n100# a_n273_131# a_n321_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 a_n129_n100# a_n177_n197# a_n225_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_63_n100# a_15_n197# a_n33_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
C0 a_159_n100# a_351_n100# 0.11fF
C1 a_n129_n100# a_n321_n100# 0.11fF
C2 a_15_n197# a_63_n100# 0.01fF
C3 a_207_n197# a_n177_n197# 0.02fF
C4 a_n81_131# a_15_n197# 0.02fF
C5 a_159_n100# a_111_131# 0.01fF
C6 a_159_n100# a_n225_n100# 0.05fF
C7 a_63_n100# a_n321_n100# 0.05fF
C8 a_303_131# a_15_n197# 0.00fF
C9 a_63_n100# a_n129_n100# 0.11fF
C10 a_207_n197# a_15_n197# 0.04fF
C11 w_n449_n200# a_n321_n100# 0.00fF
C12 w_n449_n200# a_n129_n100# 0.00fF
C13 a_n81_131# a_n129_n100# 0.01fF
C14 a_255_n100# a_n129_n100# 0.05fF
C15 a_n273_131# a_n369_n197# 0.02fF
C16 a_n369_n197# a_n177_n197# 0.04fF
C17 a_15_n197# a_n33_n100# 0.01fF
C18 a_n413_n100# a_n321_n100# 0.29fF
C19 a_n413_n100# a_n129_n100# 0.06fF
C20 w_n449_n200# a_63_n100# 0.00fF
C21 a_255_n100# a_63_n100# 0.11fF
C22 a_n33_n100# a_n321_n100# 0.06fF
C23 a_n33_n100# a_n129_n100# 0.29fF
C24 a_15_n197# a_n369_n197# 0.02fF
C25 a_255_n100# w_n449_n200# 0.00fF
C26 a_303_131# a_n81_131# 0.02fF
C27 a_207_n197# a_n81_131# 0.00fF
C28 a_303_131# a_255_n100# 0.01fF
C29 w_n449_n200# a_n413_n100# 0.00fF
C30 a_n321_n100# a_n369_n197# 0.01fF
C31 a_255_n100# a_207_n197# 0.01fF
C32 a_63_n100# a_n33_n100# 0.29fF
C33 a_303_131# a_207_n197# 0.02fF
C34 w_n449_n200# a_n33_n100# 0.00fF
C35 a_n81_131# a_n33_n100# 0.01fF
C36 a_255_n100# a_n33_n100# 0.06fF
C37 a_111_131# a_n273_131# 0.02fF
C38 a_n273_131# a_n225_n100# 0.01fF
C39 a_111_131# a_n177_n197# 0.00fF
C40 a_159_n100# a_n129_n100# 0.06fF
C41 a_n225_n100# a_n177_n197# 0.01fF
C42 a_n81_131# a_n369_n197# 0.00fF
C43 a_n413_n100# a_n33_n100# 0.05fF
C44 a_111_131# a_15_n197# 0.02fF
C45 a_159_n100# a_63_n100# 0.29fF
C46 a_n413_n100# a_n369_n197# 0.01fF
C47 a_159_n100# w_n449_n200# 0.00fF
C48 a_255_n100# a_159_n100# 0.29fF
C49 a_63_n100# a_351_n100# 0.06fF
C50 a_n273_131# a_n177_n197# 0.02fF
C51 a_n225_n100# a_n321_n100# 0.29fF
C52 a_n129_n100# a_n225_n100# 0.29fF
C53 w_n449_n200# a_351_n100# 0.00fF
C54 a_207_n197# a_159_n100# 0.01fF
C55 a_255_n100# a_351_n100# 0.29fF
C56 a_303_131# a_351_n100# 0.01fF
C57 a_159_n100# a_n33_n100# 0.11fF
C58 a_111_131# a_63_n100# 0.01fF
C59 a_15_n197# a_n273_131# 0.00fF
C60 a_63_n100# a_n225_n100# 0.06fF
C61 a_n81_131# a_111_131# 0.04fF
C62 a_15_n197# a_n177_n197# 0.04fF
C63 w_n449_n200# a_n225_n100# 0.00fF
C64 a_n33_n100# a_351_n100# 0.05fF
C65 a_303_131# a_111_131# 0.04fF
C66 a_n273_131# a_n321_n100# 0.01fF
C67 a_207_n197# a_111_131# 0.02fF
C68 a_n129_n100# a_n177_n197# 0.01fF
C69 a_n413_n100# a_n225_n100# 0.11fF
C70 a_n33_n100# a_n225_n100# 0.11fF
C71 a_n81_131# a_n273_131# 0.04fF
C72 a_n81_131# a_n177_n197# 0.02fF
C73 a_351_n100# VSUBS 0.03fF
C74 a_255_n100# VSUBS 0.03fF
C75 a_159_n100# VSUBS 0.03fF
C76 a_63_n100# VSUBS 0.03fF
C77 a_n33_n100# VSUBS 0.03fF
C78 a_n129_n100# VSUBS 0.03fF
C79 a_n225_n100# VSUBS 0.03fF
C80 a_n321_n100# VSUBS 0.03fF
C81 a_n413_n100# VSUBS 0.03fF
C82 a_207_n197# VSUBS 0.12fF
C83 a_15_n197# VSUBS 0.12fF
C84 a_n177_n197# VSUBS 0.12fF
C85 a_n369_n197# VSUBS 0.12fF
C86 a_303_131# VSUBS 0.12fF
C87 a_111_131# VSUBS 0.12fF
C88 a_n81_131# VSUBS 0.12fF
C89 a_n273_131# VSUBS 0.12fF
C90 w_n449_n200# VSUBS 1.06fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DM32AP VSUBS a_15_n100# a_n33_n188# a_n73_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
C0 a_15_n100# a_n73_n100# 0.34fF
C1 a_n33_n188# a_n73_n100# 0.03fF
C2 a_15_n100# a_n33_n188# 0.03fF
C3 a_15_n100# VSUBS 0.03fF
C4 a_n73_n100# VSUBS 0.03fF
C5 a_n33_n188# VSUBS 0.19fF
.ends

.subckt sky130_fd_pr__pfet_01v8_CW6TWB VSUBS a_n33_n197# w_n109_n200# a_15_n100# a_n73_n100#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n109_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
C0 a_15_n100# a_n33_n197# 0.03fF
C1 a_n73_n100# a_15_n100# 0.34fF
C2 w_n109_n200# a_n73_n100# 0.00fF
C3 w_n109_n200# a_15_n100# 0.00fF
C4 a_n73_n100# a_n33_n197# 0.03fF
C5 a_15_n100# VSUBS 0.03fF
C6 a_n73_n100# VSUBS 0.03fF
C7 a_n33_n197# VSUBS 0.20fF
C8 w_n109_n200# VSUBS 0.26fF
.ends

.subckt test_inverter_adj w_520_540# in sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS m1_680_300#
+ ctrl out
Xsky130_fd_pr__nfet_01v8_DM32AP_0 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS
+ in out sky130_fd_pr__nfet_01v8_DM32AP
Xsky130_fd_pr__pfet_01v8_CW6TWB_0 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS in w_520_540#
+ m1_680_300# out sky130_fd_pr__pfet_01v8_CW6TWB
Xsky130_fd_pr__pfet_01v8_CW6TWB_1 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS ctrl w_520_540#
+ w_520_540# m1_680_300# sky130_fd_pr__pfet_01v8_CW6TWB
C0 in m1_680_300# 0.27fF
C1 m1_680_300# ctrl 0.26fF
C2 m1_680_300# w_520_540# 0.08fF
C3 out m1_680_300# 0.07fF
C4 in ctrl 0.21fF
C5 in w_520_540# 0.04fF
C6 ctrl w_520_540# 0.47fF
C7 out in 0.78fF
C8 out ctrl 0.01fF
C9 out w_520_540# 0.06fF
C10 w_520_540# sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS 0.75fF
C11 ctrl sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS 0.14fF
C12 m1_680_300# sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS 0.12fF
C13 out sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS 0.20fF
C14 in sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS 0.68fF
.ends

.subckt test_osc_adj vdd vss ctrl0 ctrl1 out
Xsky130_fd_pr__pfet_01v8_RX8GT8_0 vss out vdd test_inverter_adj_2/in test_inverter_adj_2/in
+ test_inverter_adj_2/in vdd out vdd test_inverter_adj_2/in out sky130_fd_pr__pfet_01v8_RX8GT8
Xsky130_fd_pr__nfet_01v8_PE32AP_0 vss vdd vdd vss vdd vss ctrl0 vss test_inverter_adj_2/ctrl
+ ctrl1 test_inverter_adj_2/ctrl ctrl1 vss vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ sky130_fd_pr__nfet_01v8_PE32AP
Xsky130_fd_pr__nfet_01v8_CG72G3_0 vss out vss test_inverter_adj_2/in vss test_inverter_adj_2/in
+ sky130_fd_pr__nfet_01v8_CG72G3
Xsky130_fd_pr__pfet_01v8_RXQGT8_0 vss vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd
+ test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd
+ vdd sky130_fd_pr__pfet_01v8_RXQGT8
Xtest_inverter_adj_0 vdd test_inverter_adj_0/in vss test_inverter_adj_0/m1_680_300#
+ test_inverter_adj_2/ctrl test_inverter_adj_2/in test_inverter_adj
Xtest_inverter_adj_1 vdd test_inverter_adj_1/in vss test_inverter_adj_1/m1_680_300#
+ test_inverter_adj_2/ctrl test_inverter_adj_0/in test_inverter_adj
Xtest_inverter_adj_2 vdd test_inverter_adj_2/in vss test_inverter_adj_2/m1_680_300#
+ test_inverter_adj_2/ctrl test_inverter_adj_1/in test_inverter_adj
C0 test_inverter_adj_1/in test_inverter_adj_2/ctrl 0.33fF
C1 test_inverter_adj_2/in out 0.88fF
C2 test_inverter_adj_2/in ctrl0 0.01fF
C3 out vdd 1.33fF
C4 vdd ctrl0 0.05fF
C5 test_inverter_adj_0/in test_inverter_adj_2/ctrl 0.14fF
C6 ctrl1 ctrl0 0.01fF
C7 test_inverter_adj_0/m1_680_300# test_inverter_adj_0/in 0.09fF
C8 test_inverter_adj_2/in vdd 1.66fF
C9 out test_inverter_adj_2/ctrl 0.08fF
C10 test_inverter_adj_1/m1_680_300# vdd 0.33fF
C11 ctrl1 test_inverter_adj_2/in 0.03fF
C12 ctrl0 test_inverter_adj_2/ctrl 0.22fF
C13 ctrl1 vdd 0.07fF
C14 test_inverter_adj_2/m1_680_300# vdd 0.35fF
C15 test_inverter_adj_2/in test_inverter_adj_2/ctrl 0.45fF
C16 test_inverter_adj_2/in test_inverter_adj_1/in 0.15fF
C17 test_inverter_adj_1/m1_680_300# test_inverter_adj_1/in 0.09fF
C18 vdd test_inverter_adj_2/ctrl 4.86fF
C19 test_inverter_adj_1/in vdd 0.58fF
C20 ctrl1 test_inverter_adj_2/ctrl 0.39fF
C21 test_inverter_adj_0/in test_inverter_adj_2/in 0.20fF
C22 test_inverter_adj_0/in vdd 0.32fF
C23 test_inverter_adj_1/in vss 0.58fF
C24 test_inverter_adj_2/in vss 2.15fF
C25 vdd vss 5.51fF
C26 test_inverter_adj_2/ctrl vss 2.18fF
C27 test_inverter_adj_0/in vss 0.46fF
C28 out vss 1.03fF
C29 ctrl1 vss 0.27fF
C30 ctrl0 vss 0.12fF
.ends

