VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO test_osc_adj
  CLASS BLOCK ;
  FOREIGN test_osc_adj ;
  ORIGIN 0.100 0.400 ;
  SIZE 14.400 BY 5.300 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.100 2.100 14.300 4.900 ;
      LAYER li1 ;
        RECT 1.300 4.530 2.400 4.550 ;
        RECT 4.300 4.530 5.400 4.550 ;
        RECT 7.300 4.530 8.400 4.550 ;
        RECT 1.000 4.350 2.400 4.530 ;
        RECT 1.000 4.070 1.300 4.350 ;
        RECT 2.200 3.670 2.400 4.350 ;
        RECT 4.000 4.350 5.400 4.530 ;
        RECT 4.000 4.070 4.300 4.350 ;
        RECT 5.200 3.670 5.400 4.350 ;
        RECT 7.000 4.350 8.400 4.530 ;
        RECT 7.000 4.070 7.300 4.350 ;
        RECT 8.200 3.670 8.400 4.350 ;
        RECT 1.880 3.350 2.400 3.670 ;
        RECT 4.880 3.350 5.400 3.670 ;
        RECT 7.880 3.350 8.400 3.670 ;
        RECT 1.880 2.630 2.050 3.350 ;
        RECT 4.880 2.630 5.050 3.350 ;
        RECT 7.880 2.630 8.050 3.350 ;
        RECT 10.040 2.780 10.210 3.820 ;
        RECT 11.000 2.780 11.170 3.820 ;
        RECT 11.960 2.780 12.130 3.820 ;
        RECT 12.920 2.780 13.090 3.820 ;
        RECT 13.880 2.780 14.050 3.820 ;
        RECT 8.820 0.080 9.150 0.250 ;
        RECT 9.780 0.080 10.110 0.250 ;
        RECT 10.740 0.080 11.070 0.250 ;
        RECT 11.700 0.080 12.030 0.250 ;
      LAYER mcon ;
        RECT 1.880 2.710 2.050 3.590 ;
        RECT 4.880 2.710 5.050 3.590 ;
        RECT 7.880 2.710 8.050 3.590 ;
        RECT 10.040 2.860 10.210 3.740 ;
        RECT 11.000 2.860 11.170 3.740 ;
        RECT 11.960 2.860 12.130 3.740 ;
        RECT 12.920 2.860 13.090 3.740 ;
        RECT 13.880 2.860 14.050 3.740 ;
        RECT 8.900 0.080 9.070 0.250 ;
        RECT 9.860 0.080 10.030 0.250 ;
        RECT 10.820 0.080 10.990 0.250 ;
        RECT 11.780 0.080 11.950 0.250 ;
      LAYER met1 ;
        RECT 8.400 3.750 10.240 3.800 ;
        RECT 10.970 3.750 11.200 3.800 ;
        RECT 11.930 3.750 12.160 3.800 ;
        RECT 12.890 3.750 13.120 3.800 ;
        RECT 13.850 3.750 14.080 3.800 ;
        RECT 1.850 3.450 2.080 3.650 ;
        RECT 4.850 3.450 5.080 3.650 ;
        RECT 7.850 3.450 8.080 3.650 ;
        RECT 8.400 3.450 10.350 3.750 ;
        RECT 10.900 3.450 11.300 3.750 ;
        RECT 11.850 3.450 12.250 3.750 ;
        RECT 12.800 3.450 13.200 3.750 ;
        RECT 13.750 3.450 14.150 3.750 ;
        RECT 1.850 2.750 2.850 3.450 ;
        RECT 4.850 2.750 5.850 3.450 ;
        RECT 7.850 3.400 10.240 3.450 ;
        RECT 7.850 2.750 8.850 3.400 ;
        RECT 10.010 2.800 10.240 3.400 ;
        RECT 10.970 2.800 11.200 3.450 ;
        RECT 11.930 2.800 12.160 3.450 ;
        RECT 12.890 2.800 13.120 3.450 ;
        RECT 13.850 2.800 14.080 3.450 ;
        RECT 1.850 2.650 2.080 2.750 ;
        RECT 4.850 2.650 5.080 2.750 ;
        RECT 7.850 2.650 8.400 2.750 ;
        RECT 8.200 0.250 8.400 2.650 ;
        RECT 8.840 0.250 9.130 0.280 ;
        RECT 9.800 0.250 10.090 0.280 ;
        RECT 10.760 0.250 11.050 0.280 ;
        RECT 11.720 0.250 12.010 0.280 ;
        RECT 8.200 0.050 12.010 0.250 ;
      LAYER via ;
        RECT 10.000 3.450 10.300 3.750 ;
        RECT 10.950 3.450 11.250 3.750 ;
        RECT 11.900 3.450 12.200 3.750 ;
        RECT 12.850 3.450 13.150 3.750 ;
        RECT 13.800 3.450 14.100 3.750 ;
        RECT 2.200 2.750 2.800 3.450 ;
        RECT 5.200 2.750 5.800 3.450 ;
        RECT 8.200 2.750 8.800 3.450 ;
      LAYER met2 ;
        RECT 2.200 2.700 2.800 3.500 ;
        RECT 5.200 2.700 5.800 3.500 ;
        RECT 8.200 2.700 8.800 3.500 ;
        RECT 10.000 3.400 14.100 3.800 ;
      LAYER via2 ;
        RECT 2.200 2.750 2.800 3.450 ;
        RECT 5.200 2.750 5.800 3.450 ;
        RECT 8.200 2.750 8.800 3.450 ;
      LAYER met3 ;
        RECT 2.150 3.400 2.850 3.475 ;
        RECT 5.150 3.400 5.850 3.475 ;
        RECT 8.150 3.400 8.850 3.475 ;
        RECT 2.150 2.800 8.850 3.400 ;
        RECT 2.150 2.725 2.850 2.800 ;
        RECT 5.150 2.725 5.850 2.800 ;
        RECT 8.150 2.725 8.850 2.800 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 9.140 0.420 9.310 1.460 ;
        RECT 10.100 0.420 10.270 1.460 ;
        RECT 11.060 0.420 11.230 1.460 ;
        RECT 12.020 0.420 12.190 1.460 ;
      LAYER mcon ;
        RECT 9.140 0.500 9.310 1.380 ;
        RECT 10.100 0.500 10.270 1.380 ;
        RECT 11.060 0.500 11.230 1.380 ;
        RECT 12.020 0.500 12.190 1.380 ;
      LAYER met1 ;
        RECT 9.110 0.800 9.340 1.440 ;
        RECT 10.070 0.800 10.300 1.440 ;
        RECT 11.030 0.800 11.260 1.440 ;
        RECT 11.990 0.800 12.220 1.440 ;
        RECT 9.000 0.500 9.400 0.800 ;
        RECT 10.000 0.500 10.400 0.800 ;
        RECT 10.950 0.500 11.350 0.800 ;
        RECT 11.900 0.500 12.300 0.800 ;
        RECT 9.110 0.440 9.340 0.500 ;
        RECT 10.070 0.440 10.300 0.500 ;
        RECT 11.030 0.440 11.260 0.500 ;
        RECT 11.990 0.440 12.220 0.500 ;
      LAYER via ;
        RECT 9.050 0.500 9.350 0.800 ;
        RECT 10.050 0.500 10.350 0.800 ;
        RECT 11.000 0.500 11.300 0.800 ;
        RECT 11.950 0.500 12.250 0.800 ;
      LAYER met2 ;
        RECT 1.000 0.700 1.400 1.300 ;
        RECT 4.000 0.700 4.400 1.300 ;
        RECT 7.000 0.850 7.400 1.300 ;
        RECT 7.000 0.700 12.250 0.850 ;
        RECT 7.100 0.450 12.250 0.700 ;
      LAYER via2 ;
        RECT 1.000 0.750 1.400 1.250 ;
        RECT 4.000 0.750 4.400 1.250 ;
        RECT 7.000 0.750 7.400 1.250 ;
      LAYER met3 ;
        RECT 0.900 1.200 1.500 1.350 ;
        RECT 3.900 1.200 4.500 1.350 ;
        RECT 6.900 1.200 7.500 1.350 ;
        RECT 0.900 0.800 7.500 1.200 ;
        RECT 0.900 0.650 1.500 0.800 ;
        RECT 3.900 0.650 4.500 0.800 ;
        RECT 6.900 0.650 7.500 0.800 ;
    END
  END vss
  PIN ctrl0
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT 9.300 1.630 9.630 1.800 ;
      LAYER mcon ;
        RECT 9.380 1.630 9.550 1.800 ;
      LAYER met1 ;
        RECT 9.300 1.600 9.900 1.900 ;
    END
  END ctrl0
  PIN ctrl1
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 10.260 1.630 10.590 1.800 ;
        RECT 11.220 1.630 11.550 1.800 ;
      LAYER mcon ;
        RECT 10.340 1.630 10.510 1.800 ;
        RECT 11.300 1.630 11.470 1.800 ;
      LAYER met1 ;
        RECT 10.300 1.830 11.500 1.900 ;
        RECT 10.280 1.600 11.530 1.830 ;
    END
  END ctrl1
  PIN out
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER li1 ;
        RECT 6.480 3.885 6.810 4.055 ;
        RECT 0.340 2.630 0.510 3.670 ;
        RECT 6.480 2.245 6.810 2.415 ;
        RECT 6.500 1.680 6.830 1.850 ;
        RECT 0.360 0.470 0.530 1.510 ;
        RECT 6.500 0.130 6.830 0.300 ;
      LAYER mcon ;
        RECT 6.560 3.885 6.730 4.055 ;
        RECT 0.340 2.710 0.510 3.590 ;
        RECT 6.560 2.245 6.730 2.415 ;
        RECT 6.580 1.680 6.750 1.850 ;
        RECT 0.360 0.550 0.530 1.430 ;
        RECT 6.580 0.130 6.750 0.300 ;
      LAYER met1 ;
        RECT 6.450 3.850 6.850 4.150 ;
        RECT 0.310 2.850 0.540 3.650 ;
        RECT 0.100 2.650 0.540 2.850 ;
        RECT 0.100 1.500 0.300 2.650 ;
        RECT 6.450 2.150 6.850 2.450 ;
        RECT 6.500 1.950 6.800 2.150 ;
        RECT 6.450 1.650 6.850 1.950 ;
        RECT -0.100 1.490 0.500 1.500 ;
        RECT -0.100 1.250 0.560 1.490 ;
        RECT -0.100 -0.200 0.100 1.250 ;
        RECT 0.330 0.490 0.560 1.250 ;
        RECT 6.450 0.100 6.850 0.350 ;
        RECT 6.400 0.050 6.850 0.100 ;
        RECT 6.400 -0.200 6.800 0.050 ;
        RECT -0.100 -0.400 6.800 -0.200 ;
      LAYER via ;
        RECT 6.500 3.850 6.800 4.150 ;
        RECT 6.500 2.150 6.800 2.450 ;
        RECT 6.500 1.650 6.800 1.950 ;
        RECT 6.500 0.050 6.800 0.350 ;
      LAYER met2 ;
        RECT 6.500 0.000 6.800 4.200 ;
    END
  END out
  OBS
      LAYER li1 ;
        RECT 0.480 3.885 0.810 4.055 ;
        RECT 1.580 3.885 1.910 4.055 ;
        RECT 3.480 3.885 3.810 4.055 ;
        RECT 4.580 3.885 4.910 4.055 ;
        RECT 7.580 3.885 7.910 4.055 ;
        RECT 10.680 4.035 11.010 4.205 ;
        RECT 11.640 4.035 11.970 4.205 ;
        RECT 12.600 4.035 12.930 4.205 ;
        RECT 13.560 4.035 13.890 4.205 ;
        RECT 0.780 2.630 0.950 3.670 ;
        RECT 1.440 2.630 1.610 3.670 ;
        RECT 3.340 2.630 3.510 3.670 ;
        RECT 3.780 2.630 3.950 3.670 ;
        RECT 4.440 2.630 4.610 3.670 ;
        RECT 6.340 2.630 6.510 3.670 ;
        RECT 6.780 2.630 6.950 3.670 ;
        RECT 7.440 2.630 7.610 3.670 ;
        RECT 10.520 2.780 10.690 3.820 ;
        RECT 11.480 2.780 11.650 3.820 ;
        RECT 12.440 2.780 12.610 3.820 ;
        RECT 13.400 2.780 13.570 3.820 ;
        RECT 0.480 2.245 0.810 2.415 ;
        RECT 1.580 2.245 1.910 2.415 ;
        RECT 3.480 2.245 3.810 2.415 ;
        RECT 4.580 2.245 4.910 2.415 ;
        RECT 7.580 2.245 7.910 2.415 ;
        RECT 10.200 2.395 10.530 2.565 ;
        RECT 11.160 2.395 11.490 2.565 ;
        RECT 12.120 2.395 12.450 2.565 ;
        RECT 13.080 2.395 13.410 2.565 ;
        RECT 0.500 1.680 0.830 1.850 ;
        RECT 3.500 1.680 3.830 1.850 ;
        RECT 0.800 1.250 0.970 1.510 ;
        RECT 1.400 1.250 1.800 1.330 ;
        RECT 0.800 0.750 1.800 1.250 ;
        RECT 0.800 0.470 0.970 0.750 ;
        RECT 1.400 0.670 1.800 0.750 ;
        RECT 3.360 0.470 3.530 1.510 ;
        RECT 3.800 1.250 3.970 1.510 ;
        RECT 4.400 1.250 4.800 1.330 ;
        RECT 3.800 0.750 4.800 1.250 ;
        RECT 3.800 0.470 3.970 0.750 ;
        RECT 4.400 0.670 4.800 0.750 ;
        RECT 6.360 0.470 6.530 1.510 ;
        RECT 6.800 1.250 6.970 1.510 ;
        RECT 7.400 1.250 7.800 1.330 ;
        RECT 6.800 0.750 7.800 1.250 ;
        RECT 6.800 0.470 6.970 0.750 ;
        RECT 7.400 0.670 7.800 0.750 ;
        RECT 8.660 0.420 8.830 1.460 ;
        RECT 9.620 0.420 9.790 1.460 ;
        RECT 10.580 0.420 10.750 1.460 ;
        RECT 11.540 0.420 11.710 1.460 ;
        RECT 0.500 0.130 0.830 0.300 ;
        RECT 3.500 0.130 3.830 0.300 ;
      LAYER mcon ;
        RECT 0.560 3.885 0.730 4.055 ;
        RECT 1.660 3.885 1.830 4.055 ;
        RECT 3.560 3.885 3.730 4.055 ;
        RECT 4.660 3.885 4.830 4.055 ;
        RECT 7.660 3.885 7.830 4.055 ;
        RECT 10.760 4.035 10.930 4.205 ;
        RECT 11.720 4.035 11.890 4.205 ;
        RECT 12.680 4.035 12.850 4.205 ;
        RECT 13.640 4.035 13.810 4.205 ;
        RECT 0.780 2.710 0.950 3.590 ;
        RECT 1.440 2.710 1.610 3.590 ;
        RECT 3.340 2.710 3.510 3.590 ;
        RECT 3.780 2.710 3.950 3.590 ;
        RECT 4.440 2.710 4.610 3.590 ;
        RECT 6.340 2.710 6.510 3.590 ;
        RECT 6.780 2.710 6.950 3.590 ;
        RECT 7.440 2.710 7.610 3.590 ;
        RECT 10.520 2.860 10.690 3.740 ;
        RECT 11.480 2.860 11.650 3.740 ;
        RECT 12.440 2.860 12.610 3.740 ;
        RECT 13.400 2.860 13.570 3.740 ;
        RECT 0.560 2.245 0.730 2.415 ;
        RECT 1.660 2.245 1.830 2.415 ;
        RECT 3.560 2.245 3.730 2.415 ;
        RECT 4.660 2.245 4.830 2.415 ;
        RECT 7.660 2.245 7.830 2.415 ;
        RECT 10.280 2.395 10.450 2.565 ;
        RECT 11.240 2.395 11.410 2.565 ;
        RECT 12.200 2.395 12.370 2.565 ;
        RECT 13.160 2.395 13.330 2.565 ;
        RECT 0.580 1.680 0.750 1.850 ;
        RECT 3.580 1.680 3.750 1.850 ;
        RECT 0.800 0.550 0.970 1.430 ;
        RECT 3.360 0.550 3.530 1.430 ;
        RECT 3.800 0.550 3.970 1.430 ;
        RECT 6.360 0.550 6.530 1.430 ;
        RECT 6.800 0.550 6.970 1.430 ;
        RECT 8.660 0.500 8.830 1.380 ;
        RECT 9.620 0.500 9.790 1.380 ;
        RECT 10.580 0.500 10.750 1.380 ;
        RECT 11.540 0.500 11.710 1.380 ;
        RECT 0.580 0.130 0.750 0.300 ;
        RECT 3.580 0.130 3.750 0.300 ;
      LAYER met1 ;
        RECT 0.450 3.850 0.850 4.150 ;
        RECT 1.550 3.850 1.950 4.150 ;
        RECT 3.450 3.850 3.850 4.150 ;
        RECT 4.550 3.850 4.950 4.150 ;
        RECT 7.550 3.850 7.950 4.150 ;
        RECT 10.700 4.000 13.900 4.300 ;
        RECT 0.750 3.250 0.980 3.650 ;
        RECT 1.410 3.250 1.640 3.650 ;
        RECT 0.750 2.950 1.640 3.250 ;
        RECT 0.750 2.650 0.980 2.950 ;
        RECT 1.410 2.650 1.640 2.950 ;
        RECT 3.310 2.850 3.540 3.650 ;
        RECT 3.100 2.650 3.540 2.850 ;
        RECT 3.750 3.250 3.980 3.650 ;
        RECT 4.410 3.250 4.640 3.650 ;
        RECT 3.750 2.950 4.640 3.250 ;
        RECT 3.750 2.650 3.980 2.950 ;
        RECT 4.410 2.650 4.640 2.950 ;
        RECT 6.310 2.850 6.540 3.650 ;
        RECT 6.100 2.650 6.540 2.850 ;
        RECT 6.750 3.250 6.980 3.650 ;
        RECT 7.410 3.250 7.640 3.650 ;
        RECT 6.750 2.950 7.640 3.250 ;
        RECT 10.490 3.150 10.720 3.800 ;
        RECT 11.450 3.150 11.680 3.800 ;
        RECT 12.410 3.150 12.640 3.800 ;
        RECT 13.370 3.150 13.600 3.800 ;
        RECT 6.750 2.650 6.980 2.950 ;
        RECT 7.410 2.650 7.640 2.950 ;
        RECT 10.400 2.850 10.800 3.150 ;
        RECT 11.350 2.850 11.750 3.150 ;
        RECT 12.300 2.850 12.700 3.150 ;
        RECT 13.300 2.850 13.700 3.150 ;
        RECT 10.490 2.800 10.720 2.850 ;
        RECT 11.450 2.800 11.680 2.850 ;
        RECT 12.410 2.800 12.640 2.850 ;
        RECT 13.370 2.800 13.600 2.850 ;
        RECT 0.450 2.150 0.850 2.450 ;
        RECT 1.550 2.150 1.950 2.450 ;
        RECT 0.500 2.000 0.800 2.150 ;
        RECT 3.100 2.000 3.300 2.650 ;
        RECT 3.450 2.150 3.850 2.450 ;
        RECT 4.550 2.150 4.950 2.450 ;
        RECT 0.500 1.950 3.300 2.000 ;
        RECT 3.500 2.000 3.800 2.150 ;
        RECT 6.100 2.000 6.300 2.650 ;
        RECT 10.500 2.600 10.700 2.800 ;
        RECT 13.400 2.600 13.600 2.800 ;
        RECT 7.550 2.150 7.950 2.450 ;
        RECT 10.200 2.300 13.600 2.600 ;
        RECT 3.500 1.950 6.300 2.000 ;
        RECT 0.450 1.700 3.300 1.950 ;
        RECT 0.450 1.650 0.850 1.700 ;
        RECT 3.100 1.500 3.300 1.700 ;
        RECT 3.450 1.700 6.300 1.950 ;
        RECT 3.450 1.650 3.850 1.700 ;
        RECT 6.100 1.500 6.300 1.700 ;
        RECT 3.100 1.490 3.500 1.500 ;
        RECT 6.100 1.490 6.500 1.500 ;
        RECT 0.770 1.250 1.000 1.490 ;
        RECT 3.100 1.250 3.560 1.490 ;
        RECT 0.770 0.750 1.400 1.250 ;
        RECT 0.770 0.490 1.000 0.750 ;
        RECT 3.330 0.490 3.560 1.250 ;
        RECT 3.770 1.250 4.000 1.490 ;
        RECT 6.100 1.250 6.560 1.490 ;
        RECT 3.770 0.750 4.400 1.250 ;
        RECT 3.770 0.490 4.000 0.750 ;
        RECT 6.330 0.490 6.560 1.250 ;
        RECT 6.770 1.250 7.000 1.490 ;
        RECT 8.630 1.400 8.860 1.440 ;
        RECT 9.590 1.400 9.820 1.440 ;
        RECT 10.550 1.400 10.780 1.440 ;
        RECT 11.510 1.400 11.740 1.440 ;
        RECT 6.770 0.750 7.400 1.250 ;
        RECT 8.550 1.100 8.950 1.400 ;
        RECT 9.500 1.100 9.900 1.400 ;
        RECT 10.450 1.100 10.850 1.400 ;
        RECT 11.450 1.100 11.850 1.400 ;
        RECT 6.770 0.490 7.000 0.750 ;
        RECT 8.630 0.440 8.860 1.100 ;
        RECT 9.590 0.440 9.820 1.100 ;
        RECT 10.550 0.440 10.780 1.100 ;
        RECT 11.510 0.440 11.740 1.100 ;
        RECT 0.450 0.050 0.850 0.350 ;
        RECT 3.450 0.050 3.850 0.350 ;
      LAYER via ;
        RECT 0.500 3.850 0.800 4.150 ;
        RECT 1.600 3.850 1.900 4.150 ;
        RECT 3.500 3.850 3.800 4.150 ;
        RECT 4.600 3.850 4.900 4.150 ;
        RECT 7.600 3.850 7.900 4.150 ;
        RECT 10.450 2.850 10.750 3.150 ;
        RECT 11.400 2.850 11.700 3.150 ;
        RECT 12.350 2.850 12.650 3.150 ;
        RECT 13.350 2.850 13.650 3.150 ;
        RECT 0.500 2.150 0.800 2.450 ;
        RECT 1.600 2.150 1.900 2.450 ;
        RECT 3.500 2.150 3.800 2.450 ;
        RECT 4.600 2.150 4.900 2.450 ;
        RECT 7.600 2.150 7.900 2.450 ;
        RECT 0.500 1.650 0.800 1.950 ;
        RECT 3.500 1.650 3.800 1.950 ;
        RECT 8.600 1.100 8.900 1.400 ;
        RECT 9.550 1.100 9.850 1.400 ;
        RECT 10.500 1.100 10.800 1.400 ;
        RECT 11.500 1.100 11.800 1.400 ;
        RECT 0.500 0.050 0.800 0.350 ;
        RECT 3.500 0.050 3.800 0.350 ;
      LAYER met2 ;
        RECT 1.600 4.400 9.400 4.700 ;
        RECT 0.500 0.000 0.800 4.200 ;
        RECT 1.600 2.100 1.900 4.400 ;
        RECT 3.500 0.000 3.800 4.200 ;
        RECT 4.600 2.100 4.900 4.400 ;
        RECT 7.600 2.100 7.900 4.400 ;
        RECT 9.100 3.200 9.400 4.400 ;
        RECT 9.100 3.150 10.750 3.200 ;
        RECT 11.400 3.150 11.700 3.200 ;
        RECT 12.350 3.150 12.650 3.200 ;
        RECT 13.350 3.150 13.650 3.200 ;
        RECT 9.100 2.800 13.700 3.150 ;
        RECT 9.100 1.450 9.400 2.800 ;
        RECT 8.600 1.050 11.800 1.450 ;
  END
END test_osc_adj
END LIBRARY

