* NGSPICE file created from test_osc_adj.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_RX8GT8 VSUBS a_n33_n100# w_n257_n200# a_n177_n197#
+ a_n81_131# a_15_n197# a_63_n100# a_n221_n100# a_n129_n100# a_111_131# a_159_n100#
X0 a_159_n100# a_111_131# a_63_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_n33_n100# a_n81_131# a_n129_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_n129_n100# a_n177_n197# a_n221_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 a_63_n100# a_15_n197# a_n33_n100# w_n257_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PE32AP VSUBS a_63_n188# a_n129_n188# a_n81_n100# a_255_n188#
+ a_n273_n100# a_n225_122# a_111_n100# a_n177_n100# a_n33_122# a_15_n100# a_159_122#
+ a_303_n100# a_n321_n188# a_207_n100# a_n365_n100#
X0 a_15_n100# a_n33_122# a_n81_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X1 a_n273_n100# a_n321_n188# a_n365_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X2 a_n177_n100# a_n225_122# a_n273_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X3 a_303_n100# a_255_n188# a_207_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X4 a_207_n100# a_159_122# a_111_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X5 a_n81_n100# a_n129_n188# a_n177_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X6 a_111_n100# a_63_n188# a_15_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_CG72G3 VSUBS a_n33_n100# a_63_n100# a_n81_n188# a_n125_n100#
+ a_15_122#
X0 a_63_n100# a_15_122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n188# a_n125_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_RXQGT8 VSUBS a_n33_n100# a_n321_n100# a_n273_131#
+ a_n177_n197# a_n81_131# a_15_n197# a_n225_n100# w_n449_n200# a_63_n100# a_n129_n100#
+ a_303_131# a_n369_n197# a_351_n100# a_207_n197# a_255_n100# a_111_131# a_n413_n100#
+ a_159_n100#
X0 a_351_n100# a_303_131# a_255_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_255_n100# a_207_n197# a_159_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_159_n100# a_111_131# a_63_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 a_n33_n100# a_n81_131# a_n129_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 a_n321_n100# a_n369_n197# a_n413_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_n225_n100# a_n273_131# a_n321_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 a_n129_n100# a_n177_n197# a_n225_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_63_n100# a_15_n197# a_n33_n100# w_n449_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_DM32AP VSUBS a_15_n100# a_n33_n188# a_n73_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_CW6TWB VSUBS a_n33_n197# w_n109_n200# a_15_n100# a_n73_n100#
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n109_n200# sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends

.subckt test_inverter_adj w_520_540# in sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS ctrl
+ out
Xsky130_fd_pr__nfet_01v8_DM32AP_0 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS
+ in out sky130_fd_pr__nfet_01v8_DM32AP
Xsky130_fd_pr__pfet_01v8_CW6TWB_0 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS in w_520_540#
+ m1_680_300# out sky130_fd_pr__pfet_01v8_CW6TWB
Xsky130_fd_pr__pfet_01v8_CW6TWB_1 sky130_fd_pr__pfet_01v8_CW6TWB_1/VSUBS ctrl w_520_540#
+ w_520_540# m1_680_300# sky130_fd_pr__pfet_01v8_CW6TWB
.ends

.subckt test_osc_adj vdd vss ctrl0 ctrl1 out
Xsky130_fd_pr__pfet_01v8_RX8GT8_0 vss out vdd test_inverter_adj_2/in test_inverter_adj_2/in
+ test_inverter_adj_2/in vdd out vdd test_inverter_adj_2/in out sky130_fd_pr__pfet_01v8_RX8GT8
Xsky130_fd_pr__nfet_01v8_PE32AP_0 vss vdd vdd vss vdd vss ctrl0 vss test_inverter_adj_2/ctrl
+ ctrl1 test_inverter_adj_2/ctrl ctrl1 vss vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ sky130_fd_pr__nfet_01v8_PE32AP
Xsky130_fd_pr__nfet_01v8_CG72G3_0 vss out vss test_inverter_adj_2/in vss test_inverter_adj_2/in
+ sky130_fd_pr__nfet_01v8_CG72G3
Xsky130_fd_pr__pfet_01v8_RXQGT8_0 vss vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd vdd
+ test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl
+ vdd test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl test_inverter_adj_2/ctrl vdd
+ vdd sky130_fd_pr__pfet_01v8_RXQGT8
Xtest_inverter_adj_0 vdd test_inverter_adj_0/in vss test_inverter_adj_2/ctrl test_inverter_adj_2/in
+ test_inverter_adj
Xtest_inverter_adj_1 vdd test_inverter_adj_1/in vss test_inverter_adj_2/ctrl test_inverter_adj_0/in
+ test_inverter_adj
Xtest_inverter_adj_2 vdd test_inverter_adj_2/in vss test_inverter_adj_2/ctrl test_inverter_adj_1/in
+ test_inverter_adj
.ends

